module engine_0(out,clk,sod,en, in_0_0, in_0_1, in_0_2, in_0_3, in_0_4, in_0_5, in_0_6, in_0_7, in_0_8, in_0_9, in_0_10, in_0_11, in_0_12, in_0_13);
//pcre: /A°d°v°a°n°c°e°d°\s+°S°p°y°\s+°R°e°p°o°r°t°\s+°f°o°r/smi
//block char: A[0], d[1], v[2], n[3], c[4], e[5], \x20[6], S[7], p[8], y[9], R[10], o[11], t[12], f[13], 

	input clk,sod,en;

	input in_0_0, in_0_1, in_0_2, in_0_3, in_0_4, in_0_5, in_0_6, in_0_7, in_0_8, in_0_9, in_0_10, in_0_11, in_0_12, in_0_13;
	output out;


	state_0_0 St_0 (y1,1'b0,clk,en,sod);
	assign w0 = ~y1;
	state_0_1 BS_0_1 (w1,in_0_0,clk,en,sod,w0);
	state_0_2 BS_0_2 (w2,in_0_1,clk,en,sod,w1);
	state_0_3 BS_0_3 (w3,in_0_2,clk,en,sod,w2);
	state_0_4 BS_0_4 (w4,in_0_0,clk,en,sod,w3);
	state_0_5 BS_0_5 (w5,in_0_3,clk,en,sod,w4);
	state_0_6 BS_0_6 (w6,in_0_4,clk,en,sod,w5);
	state_0_7 BS_0_7 (w7,in_0_5,clk,en,sod,w6);
	state_0_8 BS_0_8 (w8,in_0_1,clk,en,sod,w7);
	state_0_9 BS_0_9 (w9,in_0_6,clk,en,sod,w9,w8);
	state_0_10 BS_0_10 (w10,in_0_7,clk,en,sod,w9);
	state_0_11 BS_0_11 (w11,in_0_8,clk,en,sod,w10);
	state_0_12 BS_0_12 (w12,in_0_9,clk,en,sod,w11);
	state_0_13 BS_0_13 (w13,in_0_6,clk,en,sod,w13,w12);
	state_0_14 BS_0_14 (w14,in_0_10,clk,en,sod,w13);
	state_0_15 BS_0_15 (w15,in_0_5,clk,en,sod,w14);
	state_0_16 BS_0_16 (w16,in_0_8,clk,en,sod,w15);
	state_0_17 BS_0_17 (w17,in_0_11,clk,en,sod,w16);
	state_0_18 BS_0_18 (w18,in_0_10,clk,en,sod,w17);
	state_0_19 BS_0_19 (w19,in_0_12,clk,en,sod,w18);
	state_0_20 BS_0_20 (w20,in_0_6,clk,en,sod,w20,w19);
	state_0_21 BS_0_21 (w21,in_0_13,clk,en,sod,w20);
	state_0_22 BS_0_22 (w22,in_0_11,clk,en,sod,w21);
	state_0_23 BS_0_23 (w23,in_0_10,clk,en,sod,w22);
	state_0_24 BS_0_24 (out,clk,en,sod,w23);
endmodule

module state_0_0(out1,in1,clk,en,rst);
	input in1,clk,rst,en;
	output out1;
	myDff Dff (out1,in1,clk,en,rst);
endmodule

module state_0_1(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_2(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_3(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_4(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_5(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_6(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_7(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_8(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_9(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_10(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_11(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_12(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_13(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_14(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_15(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_16(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_17(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_18(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_19(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_20(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_21(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_22(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_23(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	myDff Dff (out1,w2,clk,en,rst);
endmodule

module state_0_24(out1,clk,en,rst,in0);
	input clk,rst,en,in0;
	output out1;
	wire w1;
	or(w1,out1,in0);
	myDff Dff (out1,w1,clk,en,rst);
endmodule

